module cpu
(
	input clk
);


cpu_datapath LC3b_Datapath
(
		.clk(clk)
);

endmodule : cpu