import lc3b_types::*;

module memory_module
();


endmodule : memory_module