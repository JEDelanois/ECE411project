module instruction_fetch
();


endmodule : instruction_fetch