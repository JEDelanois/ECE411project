module instruction_decode
();


endmodule : instruction_decode