import lc3b_types::*;

module cpu_control
(
		input clk
);

endmodule : cpu_control