module latch_ex_mem
(
	input clk
);



endmodule : latch_ex_mem