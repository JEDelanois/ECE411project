module latch_if_id
(
	input clk
);


endmodule : latch_if_id