import lc3b_types::*;

module DivMultUnit 
(
input clk,
input [15:0] sr1, sr2,
input lc3b_aluop aluop,


output logic [15:0] solution,
output logic stall_X
);

always_comb
begin

end


endmodule : DivMultUnit