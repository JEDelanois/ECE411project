import lc3b_types::*;

module latch_id_ex
(
	input clk
);



endmodule : latch_id_ex