import lc3b_types::*;

module instruction_decode
();


endmodule : instruction_decode