module writeback_module
();


endmodule : writeback_module