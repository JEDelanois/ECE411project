import lc3b_types::*;

module writeback_module
();


endmodule : writeback_module