module memory_module
();


endmodule : memory_module