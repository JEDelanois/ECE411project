import lc3b_types::*;

module instruction_decode
(
		input clk,
		input lc3b_control control_word,
);



endmodule : instruction_decode