import lc3b_types::*;

module execution_module
();


endmodule : execution_module