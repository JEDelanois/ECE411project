import lc3b_types::*;

module cache
(
		input clk /*,
		input pmem_resp,
		input [127:0] pmem_rdata,
		output pmem_read, pmem_write,
		output [15:0] pmem_address,
		output [127:0] pmem_wdata
		*/
);

endmodule : cache