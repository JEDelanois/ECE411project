import lc3b_types::*;

module instruction_fetch
();


endmodule : instruction_fetch