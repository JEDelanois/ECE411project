module cpu_control
(
		input clk
);

endmodule : cpu_control