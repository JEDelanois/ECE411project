import lc3b_types::*;

module latch_wb
(
	input clk
);



endmodule : latch_wb