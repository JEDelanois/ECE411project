import lc3b_types::*;

module gen_control
(
		input logic [3:0] opcode,
		output lc3b_control control_word
);

endmodule : gen_control