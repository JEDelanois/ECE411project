module execution_module
();


endmodule : execution_module