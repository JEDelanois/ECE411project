import lc3b_types::*;

module latch_ex_mem
(
	input clk
);



endmodule : latch_ex_mem