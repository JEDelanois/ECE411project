module latch_wb
(
	input clk
);



endmodule : latch_wb